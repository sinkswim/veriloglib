module device(input x, input y, output z);
endmodule;
