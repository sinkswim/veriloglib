module and2(input x, input y, output z);
	and(z, x, y);
endmodule;
