// Pulse Width Modulation peripheral
// Given the input clock it generates 8 different PWM waves on the uio output pins
// Design decisions to take:
// 1) Are duty cycles fixed or can they be selected by the user using the dip switch?

module pwm
#()
();
endmodule